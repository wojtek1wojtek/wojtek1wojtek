   lsilogic           >� g�   vmware:key/list/(pair/(null/%3cVMWARE%2dEMPTYSTRING%3e,HMAC%2dSHA%2d1,mjY3iQOqugl1K4x2G7QCO7epbcOaNUmLKZBvPDN65Du3%2f9Si%2bYCEM3Wk3Y8k8t6E38w18KlTd9BDZIQ55Mxv2IcjGd4EIasumeuQj4a1VOmXoomY0T7YK5AHMr0xjKMqwQZWKlHxsiLLIigRdnN9Gz4EDTA%3d)) D  ��H*�r6,�$��J����E����F�J���W��ՠi`��s�pu��p�@�.��X�7F��l�%v��J�Ѵ\�Ix�V6�V)��1���a_������?v���4�Sr7�]֩�/�;Q��g�
���M��	[XI���G�~&Kld�1=�	j!�?K� 7�¹̑u��*�g�R��e���x�/�G�Ƅ9�P]vTi)�s�"WTy�P��M�����������+��Ù҃�H��!�a�V�hU�k�T�"K��i�2F��EZ��"3_����@Q�ÚҒG-�l,�p�ꜯ���=��M^�;$%>�E8Z�3�x����so���gq_��\|����X��w�Lg�Ɗt� ;q�P�\h�[o\���b#|��s�ִ}�I�D\���M�T������B�c��� Yp3�|���Q"��E��0l���C��`�̮v��<�"P��$��b��ߕۋ�7�~��mud���T�0�0]��}�ʀ�^��X��-�.t<*���q����<3�g:��	hGp�z	>����4�S�O\�� ���� ���o�{��I>�����n\� �}J6�(�9FŎ�"�ХC�����8f�9t`,�ٗ(4�xo���̿B��)��{/^�T���E���y̢,�Qjm��������Nn�p������~�u�#�"/TAc\�g������4�%}iN�����an<���DV��@߄��!]�v�e���Kei]N��|�pD4{�~���/�7��]�ǘv��'}3���L��L6;u� ������a�v���Ԁ_P��(�e>��U%j��]#>������<�֢f����H�����Z��¦������M0j��~'�ࠢ�>�װ��VC[XTe�D7�Z�E>7��?�������d揞�w
~�gk{��H�^��#���E��^��/����x;��.�W?fـ|Έ��p�B�&2���1�x�go�|C���.��� Z.^͂,h�Wck�=���_�0��*vQ�����[I�1��&*��۾@Cv���i��2��N�&h�4j2�¯��g�j���[�ѕ����Թ0�YB)aCR����/g�u��Zk���9����r�g-Y2/�h$�|�k�#69&��դ4�q�E�z'����Hf�ߍ�t.Ƥ��C�L:�ֱ²HUscT��=�>��#)C�/	�?J�H.Ew�Yr_���/	n�<�4'��G��f�D�q��m���6��]	Q�!c�"��$]B"hG���$�mm��4�Pp�ĕs�gm���sX�$O����=�~������ܐׅ��q�"�hYoR�.l�vI3���o���tĥ�.Vjv�m��7:&�o�Ȑ���u[��V�Piwk�U՚���M	�Zjj����e�����Ƶ��<��<mފ<JZ�LF���f!�xO�M(��Dw�|���_4a���s��F�����m�e��-�0J:	�fB�L�e̓Z�&�L��ܛT.�V�]!_��	 �k�6�g#�U[*_�q�DF(p8��U�ɃB.���h�殑V�p��l�o���i��U��